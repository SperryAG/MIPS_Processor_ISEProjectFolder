----------------------------------------------------------------------------------
-- Create Date:    18:38:32 01/16/2016 
-- Module Name:    ROM_512x32Bit - Behavioral 
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- LIBRARIES / PACKAGES
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use STD.TEXTIO.all;
use IEEE.NUMERIC_STD.all;
----------------------------------------------------------------------------------
-- ENTITY
----------------------------------------------------------------------------------
ENTITY ROM_512x32Bit IS
	PORT(
		addr   : IN    std_logic_vector(31 DOWNTO 0);
		dataIO : INOUT std_logic_vector(31 DOWNTO 0)
	);
END ROM_512x32Bit;
----------------------------------------------------------------------------------
-- ARCHITECTURE
----------------------------------------------------------------------------------
architecture Behavioral of ROM_512x32Bit is
begin
	-- pragma synthesis_off
	process is
		file mem_file: TEXT;
		variable L: line;
		variable ch: character;
		variable i, index, result: integer;
		type ramtype is array (511 downto 0) of STD_LOGIC_VECTOR(31 downto 0);
		variable mem: ramtype;
	begin
		-- initialize memory from file
		for i in 0 to 511 loop -- set all contents low
			mem(i) := (others => '0');
		end loop;

		index := 0;
		FILE_OPEN (mem_file, "memfile.dat", READ_MODE);
		while not endfile(mem_file) loop
		readline(mem_file, L);
		result := 0;

		for i in 1 to 8 loop
			read (L, ch);
			if '0' <= ch and ch <= '9' then
			result := character'pos(ch) - character'pos('0');
			elsif 'a' <= ch and ch <= 'f' then
			result := character'pos(ch) - character'pos('a')+10;
			else report "Format error on line" & integer'
			image(index) severity error;
			end if;
			mem(index)(35-i*4 downto 32-i*4) := std_logic_vector(to_unsigned(result,4));
			end loop;
			index := index + 1;
		end loop;
		-- read memory
		loop
			dataIO <= mem(to_integer(unsigned(addr(8 DOWNTO 0))));
			wait on addr;
		end loop;
	end process;
	-- pragma synthesis_on
end;